class FlyWithWings implements FlyBehavior;
   virtual function void fly();
      $display("I'm flying");
   endfunction // fly
endclass // FlyWithWings
