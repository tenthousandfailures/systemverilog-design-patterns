interface class Observer;
    pure virtual function void update(shortreal temperature, shortreal humidity, shortreal pressure);
endclass // Observer
    
