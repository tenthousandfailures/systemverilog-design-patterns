interface class QuackBehavior;
   pure virtual function void quack();
endclass // interface

