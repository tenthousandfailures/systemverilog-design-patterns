class Squeak implements QuackBehavior;
   virtual function void quack();
      $display("Squeak");
   endfunction // quack
endclass // Squeak
