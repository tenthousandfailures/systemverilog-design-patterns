class Quack implements QuackBehavior;
   virtual function void quack();
      $display("Quack");
   endfunction // quack
endclass // Quack
