virtual class CondimentDecorator extends Beverage;
	 pure virtual function string getDescription();
endclass
