interface class Observer;
   pure virtual local function void update(shortreal temperature, shortreal humidity, shortreal pressure);
   endclass // Observer

