interface class FlyBehavior;
    pure virtual function void fly();
endclass // FlyBehavior
    
