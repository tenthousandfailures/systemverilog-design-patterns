class Espresso extends Beverage;

	 function new();
      description = "Espresso";
	 endfunction

	 virtual function real cost();
      return 1.99;
	 endfunction

endclass


